`ifndef MY_DUT_SV
`define MY_DUT_SV

module my_dut(clk, rst_n, bus_cmd_valid, bus_op, bus_addr, bus_wr_data, bus_rd_data, rxd, rx_dv, txd, tx_en);
	input clk;
	input rst_n;
	input bus_cmd_valid;
	input bus_op;
	input[15:0] bus_addr;
	input[15:0] bus_wr_data;
	output[15:0] bus_rd_data;
	input[7:0] rxd;
	input rx_dv;
	output[7:0] txd;
	output tx_en;

	reg[7:0] txd;
	reg tx_en;
	reg invert;
	reg [31:0] counter;

always @(posedge clk) begin
	if(!rst_n) begin
		txd <= 8'b0;
		tx_en <= 1'b0;
	end
	else if(invert) begin
		txd <= ~rxd;
		tx_en <= rx_dv;
	end
	else begin
		txd <= rxd;
		tx_en <= rx_dv;
	end
end

always @(posedge clk) begin
	if(!rst_n) begin
		invert = 1'b0;
	end
	else if(bus_cmd_valid && bus_op) begin
		case(bus_addr)
			16'h9: begin
				invert <= bus_wr_data[0];
			end
			default: begin
			end
		endcase
	end
end

reg[15:0] bus_rd_data;
always @(posedge clk) begin
	if(!rst_n) begin
		bus_rd_data <= 0;
	end
	else if(bus_cmd_valid && (!bus_op)) begin
		case(bus_addr)
			16'h9: begin
				bus_rd_data <= {15'b0, invert};
			end
			default: begin
				bus_rd_data <= 16'b0;
			end
		endcase
	end
end

endmodule
`endif
